// Code your design here
`include "Definitions.sv"
`include "TopLevel.sv"
`include "Immediate_LUT.sv"
`include "lut.sv"
`include "Ctrl.sv"
`include "InstFetch.sv"
`include "RegFile.sv"
`include "InstROM.sv"
`include "ALU.sv"
`include "DataMem.sv"


