// Code your testbench here
// or browse Examples
`include "program1_tb.sv"